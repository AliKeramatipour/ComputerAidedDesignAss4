library verilog;
use verilog.vl_types.all;
entity TBFD is
end TBFD;
